module block_update (ClkPort, number1, number2, number3, number4, number5, number6, number7, number8, number9, 
			number10, number11, number12, number13, number14, number15, number16, x, y);

input ClkPort;

input [10:0] number1;
input [10:0] number2;
input [10:0] number3;
input [10:0] number4;
input [10:0] number5;
input [10:0] number6;
input [10:0] number7;
input [10:0] number8;
input [10:0] number9;
input [10:0] number10;
input [10:0] number11;
input [10:0] number12;
input [10:0] number13;
input [10:0] number14;
input [10:0] number15;
input [10:0] number16;

input [9:0] x;
input [9:0] y;

output [2:0] red;
output [2:0] green;
output [1:0] blue;

box box_00 (10, 12, number1, x, y);
box box_01 (175, 12, number2, x, y);
box box_02 (325, 12, number3, x, y);
box box_03 (485, 12, number4, x, y);

box box_10 (10, 129, number5, x, y);
box box_11 (175, 129, number6, x, y);
box box_12 (325, 129, number7, x, y);
box box_13 (485, 129, number8, x, y);

box box_20 (10, 246, number9, x, y);
box box_21 (175, 246, number10, x, y);
box box_22 (325, 246, number11, x, y);
box box_23 (485, 246, number12, x, y);

box box_30 (10, 363, number13, x, y);
box box_31 (175, 363, number14, x, y);
box box_32 (325, 363, number15, x, y);
box box_33 (485, 363, number16, x, y);


always @ (posedge ClkPort)
	begin 
		case (number1)
			11'b00000000000: 
				box_00 (10,12,0,x,y);
			11'b00000000001:
				box_00 (10,12,2,x,y);
			11'b00000000010:
				box_00 (10,12,4,x,y);
			11'b00000000100:
				box_00 (10,12,8,x,y);	
			11'b00000001000:
				box_00 (10,12,16,x,y);
			11'b00000010000:
				box_00 (10,12,32,x,y);
			11'b00000100000:
				box_00 (10,12,64,x,y);
			11'b00001000000:
				box_00 (10,12,128,x,y);
			11'b00010000000:
				box_00 (10,12,256,x,y);
			11'b00100000000:
				box_00 (10,12,512,x,y);
			11'b01000000000:
				box_00 (10,12,1024,x,y);
			11'b10000000000:
				box_00 (10,12,2048,x,y);
	end
	
		case (number2)
			11'b00000000000: 
				box_01 (175,12,0,x,y);
			11'b00000000001:
				box_01 (175,12,2,x,y);
			11'b00000000010:
				box_01 (175,12,4,x,y);
			11'b00000000100:
				box_01 (175,12,8,x,y);	
			11'b00000001000:
				box_01 (175,12,16,x,y);
			11'b00000010000:
				box_01 (175,12,32,x,y);
			11'b00000100000:
				box_01 (175,12,64,x,y);
			11'b00001000000:
				box_01 (175,12,128,x,y);
			11'b00010000000:
				box_01 (175,12,256,x,y);
			11'b00100000000:
				box_01 (175,12,512,x,y);
			11'b01000000000:
				box_01 (175,12,1024,x,y);
			11'b10000000000:
				box_01 (175,12,2048,x,y);
	end
	
		case (number3)
			11'b00000000000: 
				box_02 (325,12,0,x,y);
			11'b00000000001:
				box_02 (325,12,2,x,y);
			11'b00000000010:
				box_02 (325,12,4,x,y);
			11'b00000000100:
				box_02 (325,12,8,x,y);	
			11'b00000001000:
				box_02 (325,12,16,x,y);
			11'b00000010000:
				box_02 (325,12,32,x,y);
			11'b00000100000:
				box_02 (325,12,64,x,y);
			11'b00001000000:
				box_02 (325,12,128,x,y);
			11'b00010000000:
				box_02 (325,12,256,x,y);
			11'b00100000000:
				box_02 (325,12,512,x,y);
			11'b01000000000:
				box_02 (325,12,1024,x,y);
			11'b10000000000:
				box_02 (325,12,2048,x,y);
	end
	
		case (number4)
			11'b00000000000: 
				box_03 (485,12,0,x,y);
			11'b00000000001:
				box_03 (485,12,2,x,y);
			11'b00000000010:
				box_03 (485,12,4,x,y);
			11'b00000000100:
				box_03 (485,12,8,x,y);	
			11'b00000001000:
				box_03 (485,12,16,x,y);
			11'b00000010000:
				box_03 (485,12,32,x,y);
			11'b00000100000:
				box_03 (485,12,64,x,y);
			11'b00001000000:
				box_03 (485,12,128,x,y);
			11'b00010000000:
				box_03 (485,12,256,x,y);
			11'b00100000000:
				box_03 (485,12,512,x,y);
			11'b01000000000:
				box_03 (485,12,1024,x,y);
			11'b10000000000:
				box_03 (485,12,2048,x,y);
	end
	
		case (number5)
			11'b00000000000: 
				box_10 (10,129,0,x,y);
			11'b00000000001:
				box_10 (10,129,2,x,y);
			11'b00000000010:
				box_10 (10,129,4,x,y);
			11'b00000000100:
				box_10 (10,129,8,x,y);	
			11'b00000001000:
				box_10 (10,129,16,x,y);
			11'b00000010000:
				box_10 (10,129,32,x,y);
			11'b00000100000:
				box_10 (10,129,64,x,y);
			11'b00001000000:
				box_10 (10,129,128,x,y);
			11'b00010000000:
				box_10 (10,129,256,x,y);
			11'b00100000000:
				box_10 (10,129,512,x,y);
			11'b01000000000:
				box_10 (10,129,1024,x,y);
			11'b10000000000:
				box_10 (10,129,2048,x,y);
	end
		
		case (number6)
			11'b00000000000: 
				box_11 (175,129,0,x,y);
			11'b00000000001:
				box_11 (175,129,2,x,y);
			11'b00000000010:
				box_11 (175,129,4,x,y);
			11'b00000000100:
				box_11 (175,129,8,x,y);	
			11'b00000001000:
				box_11 (175,129,16,x,y);
			11'b00000010000:
				box_11 (175,129,32,x,y);
			11'b00000100000:
				box_11 (175,129,64,x,y);
			11'b00001000000:
				box_11 (175,129,128,x,y);
			11'b00010000000:
				box_11 (175,129,256,x,y);
			11'b00100000000:
				box_11 (175,129,512,x,y);
			11'b010000000000:
				box_11 (175,129,1024,x,y);
			11'b100000000000:
				box_10 (175,129,2048,x,y);
	end
	
		case (number7)
			11'b00000000000: 
				box_12 (325,129,0,x,y);
			11'b00000000001:
				box_12 (325,129,2,x,y);
			11'b00000000010:
				box_12 (325,129,4,x,y);
			11'b00000000100:
				box_12 (325,129,8,x,y);	
			11'b00000001000:
				box_12 (325,129,16,x,y);
			11'b00000010000:
				box_12 (325,129,32,x,y);
			11'b00000100000:
				box_12 (325,129,64,x,y);
			11'b00001000000:
				box_12 (325,129,128,x,y);
			11'b00010000000:
				box_12 (325,129,256,x,y);
			11'b00100000000:
				box_12 (325,129,512,x,y);
			11'b01000000000:
				box_12 (325,129,1024,x,y);
			11'b10000000000:
				box_12 (325,129,2048,x,y);
	end
	
		case (number8)
			11'b00000000000: 
				box_13 (485,129,0,x,y);
			11'b00000000001:
				box_13 (485,129,2,x,y);
			11'b00000000010:
				box_13 (485,129,4,x,y);
			11'b00000000100:
				box_13 (485,129,8,x,y);	
			11'b00000001000:
				box_13 (485,129,16,x,y);
			11'b00000010000:
				box_13 (485,129,32,x,y);
			11'b00000100000:
				box_13 (485,129,64,x,y);
			11'b00001000000:
				box_13 (485,129,128,x,y);
			11'b00010000000:
				box_13 (485,129,256,x,y);
			11'b00100000000:
				box_13 (485,129,512,x,y);
			11'b01000000000:
				box_13 (485,129,1024,x,y);
			11'b10000000000:
				box_13 (485,129,2048,x,y);
	end
	
		case (number9)
			11'b00000000000: 
				box_20 (10,246,0,x,y);
			11'b00000000001:
				box_20 (10,246,2,x,y);
			11'b00000000010:
				box_20 (10,246,4,x,y);
			11'b00000000100:
				box_20 (10,246,8,x,y);	
			11'b00000001000:
				box_20 (10,246,16,x,y);
			11'b00000010000:
				box_20 (10,246,32,x,y);
			11'b00000100000:
				box_20 (10,246,64,x,y);
			11'b00001000000:
				box_20 (10,246,128,x,y);
			11'b00010000000:
				box_20 (10,246,256,x,y);
			11'b00100000000:
				box_20 (10,246,512,x,y);
			11'b01000000000:
				box_20 (10,246,1024,x,y);
			11'b100000000000:
				box_20 (10,246,2048,x,y);
	end
		
		case (number10)
			11'b00000000000: 
				box_21 (175,246,0,x,y);
			11'b00000000001:
				box_21 (175,246,2,x,y);
			11'b00000000010:
				box_21 (175,246,4,x,y);
			11'b00000000100:
				box_21 (175,246,8,x,y);	
			11'b00000001000:
				box_21 (175,246,16,x,y);
			11'b00000010000:
				box_21 (175,246,32,x,y);
			11'b00000100000:
				box_21 (175,246,64,x,y);
			11'b00001000000:
				box_21 (175,246,128,x,y);
			11'b00010000000:
				box_21 (175,246,256,x,y);
			11'b00100000000:
				box_21 (175,246,512,x,y);
			11'b01000000000:
				box_21 (175,246,1024,x,y);
			11'b10000000000:
				box_21 (175,246,2048,x,y);
	end
	
		case (number11)
			11'b00000000000: 
				box_22 (325,246,0,x,y);
			11'b00000000001:
				box_22 (325,246,2,x,y);
			11'b00000000010:
				box_22 (325,246,4,x,y);
			11'b00000000100:
				box_22 (325,246,8,x,y);	
			11'b00000001000:
				box_22 (325,246,16,x,y);
			11'b00000010000:
				box_22 (325,246,32,x,y);
			11'b00000100000:
				box_22 (325,246,64,x,y);
			11'b00001000000:
				box_22 (325,246,128,x,y);
			11'b00010000000:
				box_22 (325,246,256,x,y);
			11'b00100000000:
				box_22 (325,246,512,x,y);
			11'b01000000000:
				box_22 (325,246,1024,x,y);
			11'b10000000000:
				box_22 (325,246,2048,x,y);
	end
	
		case (number12)
			11'b00000000000: 
				box_23 (485,246,0,x,y);
			11'b00000000001:
				box_23 (485,246,2,x,y);
			11'b00000000010:
				box_23 (485,246,4,x,y);
			11'b00000000100:
				box_23 (485,246,8,x,y);	
			11'b00000001000:
				box_23 (485,246,16,x,y);
			11'b00000010000:
				box_23 (485,246,32,x,y);
			11'b00000100000:
				box_23 (485,246,64,x,y);
			11'b00001000000:
				box_23 (485,246,128,x,y);
			11'b00010000000:
				box_23 (485,246,256,x,y);
			11'b00100000000:
				box_23 (485,246,512,x,y);
			11'b01000000000:
				box_23 (485,246,1024,x,y);
			11'b10000000000:
				box_23 (485,246,2048,x,y);
	end	
	
		case (number13)
			11'b00000000000: 
				box_30 (10,363,0,x,y);
			11'b00000000001:
				box_30 (10,363,2,x,y);
			11'b00000000010:
				box_30 (10,363,4,x,y);
			11'b00000000100:
				box_30 (10,363,8,x,y);	
			11'b00000001000:
				box_30 (10,363,16,x,y);
			11'b00000010000:
				box_30 (10,363,32,x,y);
			11'b00000100000:
				box_30 (10,363,64,x,y);
			11'b00001000000:
				box_30 (10,363,128,x,y);
			11'b00010000000:
				box_33 (10,363,256,x,y);
			11'b00100000000:
				box_33 (10,363,512,x,y);
			11'b01000000000:
				box_33 (10,363,1024,x,y);
			11'b10000000000:
				box_33 (10,363,2048,x,y);
	end	
		
		case (number14)
			11'b00000000000: 
				box_31 (175,363,0,x,y);
			11'b00000000001:
				box_31 (175,363,2,x,y);
			11'b00000000010:
				box_31 (175,363,4,x,y);
			11'b00000000100:
				box_31 (175,363,8,x,y);	
			11'b00000001000:
				box_31 (175,363,16,x,y);
			11'b00000010000:
				box_31 (175,363,32,x,y);
			11'b00000100000:
				box_31 (175,363,64,x,y);
			11'b00001000000:
				box_31 (175,363,128,x,y);
			11'b00010000000:
				box_31 (175,363,256,x,y);
			11'b00100000000:
				box_31 (175,363,512,x,y);
			11'b01000000000:
				box_31 (175,363,1024,x,y);
			11'b10000000000:
				box_31 (175,363,2048,x,y);
	end	
	
		case (number15)
			11'b00000000000: 
				box_32 (325,363,0,x,y);
			11'b00000000001:
				box_32 (325,363,2,x,y);
			11'b00000000010:
				box_32 (325,363,4,x,y);
			11'b00000000100:
				box_32 (325,363,8,x,y);	
			11'b00000001000:
				box_32 (325,363,16,x,y);
			11'b00000010000:
				box_32 (325,363,32,x,y);
			11'b00000100000:
				box_32 (325,363,64,x,y);
			11'b00001000000:
				box_32 (325,363,128,x,y);
			11'b00010000000:
				box_32 (325,363,256,x,y);
			11'b00100000000:
				box_32 (325,363,512,x,y);
			11'b01000000000:
				box_32 (325,363,1024,x,y);
			11'b10000000000:
				box_32 (325,363,2048,x,y);
	end	
		
		case (number16)
			11'b00000000000: 
				box_33 (485,363,0,x,y);
			11'b00000000001:
				box_33 (485,363,2,x,y);
			11'b00000000010:
				box_33 (485,363,4,x,y);
			11'b00000000100:
				box_33 (485,363,8,x,y);	
			11'b00000001000:
				box_33 (485,363,16,x,y);
			11'b00000010000:
				box_33 (485,363,32,x,y);
			11'b00000100000:
				box_33 (485,363,64,x,y);
			11'b00001000000:
				box_33 (485,363,128,x,y);
			11'b00010000000:
				box_33 (485,363,256,x,y);
			11'b00100000000:
				box_33 (485,363,512,x,y);
			11'b01000000000:
				box_33 (485,363,1024,x,y);
			11'b10000000000:
				box_33 (485,363,2048,x,y);
	end	
			
endmodule